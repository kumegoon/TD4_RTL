`define cycle               1000
`define cycle_duty          `cycle/2
`define max_cycle_count     150000
`timescale                  1ns/1ns

// module declare

module full_adder_tb;

//wire and reg
    reg [1:0]       IN_Y;
    reg [1:0]       IN_DATA;
    reg [1:0]       CIN;
    reg [1:0]       IN_Y;
    reg [1:0]       IN_Y;